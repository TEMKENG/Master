library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity VISCY_CPU_TB IS
end VISCY_CPU_TB;

architecture BEHAVIOR of VISCY_CPU_TB is

-- Component Declaration for the Unit
component VISCY_CPU
	port (
		clk, reset, ready : in std_logic;
		rd, wr : out std_logic;
		adr
		: out std_logic_vector (15 downto 0);
		rdata : in std_logic_vector (15 downto 0);
		wdata : out std_logic_vector (15 downto 0)
	);
end component;

-- Signals...
signal clk, reset, ready, rd, wr: std_logic;
signal adr, rdata, wdata: std_logic_vector (15 downto 0);

-- Parameters...
constant clk_period: time := 10 ns;
constant mem_delay: time := 25 ns;

 -- Memory content (generated by viscy2l) ...
  -- type t_memory is array (0 to 271) of std_logic_vector (15 downto 0);
  -- signal mem_content: t_memory := (
      -- 16#0000# => "0100000100000001",  -- 	ldil  		r1, 1
      -- 16#0001# => "0100100100000000",  -- 	ldih 		r1, 0
      -- 16#0002# => "0100011100000000",  -- 	ldil  		r7,  0x00
      -- 16#0003# => "0100111100000001",  -- 	ldih 		r7,  0x01 ; r7:=0x0100
      -- 16#0004# => "0011000011111100",  -- 	XOR			r0, r7, r7; r0:=0
      -- 16#0005# => "0101100011100000",  -- 	st			[r7], r0 ; speichern r0 in adresse r7
      -- 16#0006# => "0100000000001000",  -- 	ldil 		r0, 0x08; ; ro:= 0x08
      -- 16#0007# => "0000011111100100",  -- 	add 		r7, r7, r1;  Zieladresse erhoehen
      -- 16#0008# => "0001000000000000",  -- 	sal 		r0, r0; shift nach links
      -- 16#0009# => "0101100011100000",  -- 	st			[r7], r0; speichern von ro in der Adresse r7
      -- 16#000a# => "0101001011100000",  -- 	ld 			r2, [r7]; Laden des Wertes von der Speicheradresse r7 in r2
      -- 16#000b# => "0001100000000000",  -- 	sar 		r0, r0; shift nach rechts
      -- 16#000c# => "0000011111100100",  -- 	add 		r7, r7, r1; Zieladresse erhoehen
      -- 16#000d# => "0101100011100000",  -- 	st			[r7], r0 ; speichern von ro in der adresse r7
      -- 16#000e# => "0100000000001111",  -- 	ldil		r0, 0x0f ;
      -- 16#000f# => "0100100011110000",  -- 	ldih		r0, 0xf0; r0 :=0xf00f
      -- 16#0010# => "0100001011110000",  -- 	ldil		r2, 0xf0
      -- 16#0011# => "0100101000001111",  -- 	ldih		r2, 0x0f; r2:=0x0ff0
      -- 16#0012# => "0000100000001000",  -- 	sub			r0, r0, r2; ro:= r0-r2
      -- 16#0013# => "0000011111100100",  -- 	add 		r7, r7, r1; Zieladresse erhoehen
      -- 16#0014# => "0101100011100000",  -- 	st			[r7], r0; speichern von ro in der Adresse r7
      -- 16#0015# => "0011100001000000",  -- 	not			r0, r2 ; ro:= not r2
      -- 16#0016# => "0000011111100100",  -- 	add 		r7, r7, r1; Zieladresse erhoehen
      -- 16#0017# => "0101100011100000",  -- 	st			[r7], r0;speichern von ro in der Adresse r7
      -- 16#0018# => "0100101000000000",  -- 	ldih		r2, 0 ;
      -- 16#0019# => "0100001000000111",  -- 	ldil		r2, 7 ; r2 := 7
      -- 16#001a# => "0100101111111111",  -- 	ldih		r3, 0xFF
      -- 16#001b# => "0100001111111111",  -- 	ldil		r3, 0xFF; r3 := 0xFFFF;
      -- 16#001c# => "0010000001001100",  -- 	and			r0, r2, r3 ; r0:= r2 and r3
      -- 16#001d# => "0000011111100100",  -- 	add 		r7, r7, r1; Zieladresse erhoehen
      -- 16#001e# => "0101100011100000",  -- 	st			[r7], r0 ;speichern von ro in der Adresse r7
      -- 16#001f# => "0100000010101010",  -- 	ldil 		r0, 0xAA
      -- 16#0020# => "0100100010101010",  -- 	ldih 		r0, 0xAA ; r0:= 0xAAAA
      -- 16#0021# => "0100001001010101",  -- 	ldil		r2, 0x55
      -- 16#0022# => "0100101001010101",  -- 	ldih		r2, 0x55 ; r2:= 0x5555
      -- 16#0023# => "0010100000001000",  -- 	or			r0, r0, r2; r0 := r0 or r2
      -- 16#0024# => "0000011111100100",  -- 	add 		r7, r7, r1 ; Zieladresse erhoehen
      -- 16#0025# => "0101100011100000",  -- 	st			[r7], r0 ; speichern von ro in der Adresse r7
      -- 16#0026# => "0100001000000101",  -- 	ldil		r2, 0x05
      -- 16#0027# => "0100101000000000",  -- 	ldih		r2, 0x00 ; r2:= ox0005
      -- 16#0028# => "0011000000000000",  -- 	xor			r0, r0, r0 ; r0 := r0 xor r0
      -- 16#0029# => "0100010000110001",  -- 	ldil		r4, end & 255 ; r4:= end(Adresse)
      -- 16#002a# => "0100110000000000",  -- 	ldih		r4, end >> 8
      -- 16#002b# => "0100001100101101",  -- 	ldil		r3, loop & 255 ;r3:= loop (Sprungadresse)
      -- 16#002c# => "0100101100000000",  -- 	ldih		r3, loop >> 8
      -- 16#002d# => "1001000010001000",  -- 	jz			r2, r4; spring auf end when r2 :=0
      -- 16#002e# => "0000000000001000",  -- 	add 		r0, r0, r2; Zieladresse erhoehen
      -- 16#002f# => "0000101001000100",  -- 	sub 		r2, r2, r1;  r2:=r2-1 ; Schleifenzaehler erniedrigen
      -- 16#0030# => "1000000001100000",  -- 	jmp 		r3 ; spring nach loop
      -- 16#0031# => "0000011111100100",  -- 	add 		r7, r7, r1 ;Zieladresse erhoehen
      -- 16#0032# => "0101100011100000",  -- 	st			[r7], r0 ; speichern von ro in der Adresse r7
      -- 16#0033# => "0100001000000010",  -- 	ldil		r2, 0x02
      -- 16#0034# => "0100101000000000",  -- 	ldih		r2, 0x00 ; r2:= ox0002
      -- 16#0035# => "0011000000000000",  -- 	xor			r0, r0, r0 ; r0:=0
      -- 16#0036# => "0000000000001000",  -- 	add 		r0, r0, r2 ;r0 := r0+r2
      -- 16#0037# => "0000101001000100",  -- 	sub 		r2, r2, r1; r2:= r2+r1
      -- 16#0038# => "0100001100110110",  -- 	ldil		r3, loop1 & 255 ; r3:= loop (Sprungadresse)
      -- 16#0039# => "0100101100000000",  -- 	ldih		r3, loop1 >> 8
      -- 16#003a# => "1001100001101000",  -- 	jnz 		r2, r3 ;  spring nach loop falls r2!=0
      -- 16#003b# => "0000011111100100",  -- 	add 		r7, r7, r1 ;Zieladresse erhoehen
      -- 16#003c# => "0101100011100000",  -- 	st			[r7], r0 ; speichern von ro in der Adresse r7
      -- 16#003d# => "1000100000000000",  -- 	halt        ;prozessor anhalten
      -- 16#0100# => "0000000000000000",  -- 	.res 16
      -- 16#0101# => "0000000000000000",
      -- 16#0102# => "0000000000000000",
      -- 16#0103# => "0000000000000000",
      -- 16#0104# => "0000000000000000",
      -- 16#0105# => "0000000000000000",
      -- 16#0106# => "0000000000000000",
      -- 16#0107# => "0000000000000000",
      -- 16#0108# => "0000000000000000",
      -- 16#0109# => "0000000000000000",
      -- 16#010a# => "0000000000000000",
      -- 16#010b# => "0000000000000000",
      -- 16#010c# => "0000000000000000",
      -- 16#010d# => "0000000000000000",
      -- 16#010e# => "0000000000000000",
      -- 16#010f# => "0000000000000000",
      -- others => "UUUUUUUUUUUUUUUU"

    -- );


 type t_memory is array (0 to 258) of std_logic_vector (15 downto 0);
  signal mem_content: t_memory := (
      16#0000# => "0100011100000000",  -- 	ldil	r7, 0x00
      16#0001# => "0100111100000001",  -- 	ldih	r7, 0x01
      16#0002# => "0101000011100000",  -- 	ld	r0, [r7]
      16#0003# => "0100011100000001",  -- 	ldil	r7, 0x01
      16#0004# => "0101000111100000",  -- 	ld	r1, [r7]
      16#0005# => "0100011100101111",  -- 	ldil	r7, result & 255 ; r7 := result(Adresse)
      16#0006# => "0100111100000000",  -- 	ldih	r7, result >> 8
      16#0007# => "1001000011100000",  -- 	jz	r0, r7
      16#0008# => "1001000011100100",  -- 	jz	r1, r7
      16#0009# => "0011011011111100",  -- 	xor r6, r7, r7 ; r6:=result :=0
      16#000a# => "0100001000000000",  -- 	ldil	r2, 0x00
      16#000b# => "0100101010000000",  -- 	ldih	r2, 0x80
      16#000c# => "0100001100010000",  -- 	ldil	r3, 16
      16#000d# => "0100101100000000",  -- 	ldih	r3, 0
      16#000e# => "0100010100000001",  -- 	ldil	r5, 1 	;r5 = 1 Konstante
      16#000f# => "0100110100000000",  -- 	ldih	r5, 0
      16#0010# => "0100011100101111",  -- 	ldil	r7, result & 255 	; r7 := result(Adresse)
      16#0011# => "0100111100000000",  -- 	ldih	r7, result >> 8
      16#0012# => "1001000011101100",  -- 	jz 		r3, r7 				; zaehler == 0
      16#0013# => "0010010000101000",  -- 	and 	r4, r1, r2
      16#0014# => "0100011100011101",  -- 	ldil	r7, addi & 255 		; r7 := addi(Adresse)
      16#0015# => "0100111100000000",  -- 	ldih	r7, addi >> 8
      16#0016# => "1001100011110000",  -- 	jnz  	r4, r7				;Springt zu addi, wenn r4 != 0
      16#0017# => "0100011100100100",  -- 	ldil	r7, mul2 & 255 		; r7 := mul2(Adresse)
      16#0018# => "0100111100000000",  -- 	ldih	r7, mul2 >> 8
      16#0019# => "1001100011111000",  -- 	jnz  	r6, r7				;Springt zu mul2, wenn r6 != 0
      16#001a# => "0100011100101010",  -- 	ldil	r7, update & 255 	; r7 := update(Adresse)
      16#001b# => "0100111100000000",  -- 	ldih	r7, update >> 8
      16#001c# => "1000000011100000",  -- 	jmp		r7					;Springt zu update
      16#001d# => "0100011100101000",  -- 	ldil	r7, muladd & 255 	; r7 := muladd(Adresse)
      16#001e# => "0100111100000000",  -- 	ldih	r7, muladd >> 8
      16#001f# => "1001100011111000",  -- 	jnz		r6, r7				;Springt zu muladd, wenn r6 != 0
      16#0020# => "0000011011000000",  -- 	add  	r6, r6, r0			;Erste Schleife Durchlauf
      16#0021# => "0100011100101010",  -- 	ldil	r7, update & 255 	; r7 := update(Adresse)
      16#0022# => "0100111100000000",  -- 	ldih	r7, update >> 8
      16#0023# => "1000000011100000",  -- 	jmp   	r7					;Springt zu update
      16#0024# => "0001011011000000",  -- 	sal r6, r6 					; r6 *=2
      16#0025# => "0100011100101010",  -- 	ldil	r7, update & 255 	; r7 := update(Adresse)
      16#0026# => "0100111100000000",  -- 	ldih	r7, update >> 8
      16#0027# => "1000000011100000",  -- 	jmp   	r7 					;Springt zu update
      16#0028# => "0001011011000000",  -- 	sal 	r6, r6 				; r6 *=2
      16#0029# => "0000011011000000",  -- 	add		r6, r6, r0			; r6 = r6 + r0 = r6 + a
      16#002a# => "0000101101110100",  -- 	sub 	r3, r3, r5 			; zaehler dekrementieren r3 -=1
      16#002b# => "0001000100100000",  -- 	sal 	r1, r1	   			; b=r1=r1*2 = b*2
      16#002c# => "0100011100010000",  -- 	ldil	r7, loop & 255 		; r7 := loop(Sprungdresse)
      16#002d# => "0100111100000000",  -- 	ldih	r7, loop >> 8
      16#002e# => "1000000011100000",  -- 	jmp		r7					;Springt zu loop
      16#002f# => "0100011100000010",  -- 	ldil	r7, 0x02 			; r7 := Ergebnis Adresse
      16#0030# => "0100111100000001",  -- 	ldih	r7, 0x01
      16#0031# => "0101100011111000",  -- 	st	[r7], r6 				; Ergebnis speichern
      16#0032# => "1000100000000000",  -- 	halt
      16#0100# => "0000000010110000",  -- .data 176, 176 					;a=(Wert=40 Adresse=0x0100) , b=(Wert=2 Adresse=0x0101)
      16#0101# => "0000000010100111",
      16#0102# => "0000000000000000", -- .res 1
      others => "UUUUUUUUUUUUUUUU"
    );



    
begin
-- Instantiate the Unit Under Test (UUT)
UUT: VISCY_CPU port map (
	clk => clk, reset => reset,
	rd => rd, wr => wr, ready => ready,
	adr => adr, rdata => rdata, wdata => wdata
);
-- Process to simulate the memory behavior...
memory : process
begin
	ready <= '0';
	wait on rd, wr;
		if rd = '1' then
			wait for mem_delay;
			if is_x (adr) then
				rdata <= (others => 'X');
			else
				rdata <= mem_content (to_integer (unsigned (adr)));
			end if;
			ready <= '1';
			wait until rd = '0';
				rdata <= (others => 'X');
			wait for mem_delay;
				ready <= '0';
		elsif wr = '1' then
			wait for mem_delay;
			if not is_x(adr) then
				mem_content (to_integer (unsigned (adr))) <= wdata;
			end if;
			ready <= '1';
			wait until wr = '0';
			wait for mem_delay;
			ready <= '0';
		end if;
end process;

-- Main testbench process...
tb : process
	procedure run_cycle is
	begin
	clk <= '0';
	wait for clk_period / 2;
	clk <= '1';
	wait for clk_period / 2;
	end procedure;
	variable nb_takt: integer :=0;
	begin
	-- SINNVOLLES HAUPTPROGRAMM UEBERLEGEN
		
	reset <= '1';
	run_cycle;
	reset <= '0';

	while nb_takt <= 10 loop
		if(rd = '0') then
			nb_takt := nb_takt + 1;
		else
			nb_takt := 0;
		end if;
		run_cycle;
			report "TEST " & integer'image(to_integer(unsigned(adr)));

	end loop;
	wait;
	-- wait forever (stop simulation)
end process;
end;

