library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity VISCY_CPU_TB IS
end VISCY_CPU_TB;

architecture BEHAVIOR of VISCY_CPU_TB is

-- Component Declaration for the Unit
component VISCY_CPU
	port (
		clk, reset, ready : in std_logic;
		rd, wr : out std_logic;
		adr
		: out std_logic_vector (15 downto 0);
		rdata : in std_logic_vector (15 downto 0);
		wdata : out std_logic_vector (15 downto 0)
	);
end component;

-- Signals...
signal clk, reset, ready, rd, wr: std_logic;
signal adr, rdata, wdata: std_logic_vector (15 downto 0);

-- Parameters...
constant clk_period: time := 10 ns;
constant mem_delay: time := 25 ns;

-- Memory content (generated by viscy2l) ...
type t_memory is array (0 to 19) of std_logic_vector (15 downto 0);
  signal mem_content: t_memory := (
      16#0000# => "0011000000000000",  -- 			XOR r0, r0, r0	; r0 beinhaltet nur '0'
      16#0001# => "0100100000000001",  -- 			LDIH r0, 0x01  	; r0 := 0x100
      16#0002# => "0101000100000000",  -- 			LD r1, [r0]   	; 1. Wert in r1
      16#0003# => "0011000000000000",  -- 			XOR   r0, r0, r0
      16#0004# => "0100000000000001",  -- 			LDIL  r0, 0x01
      16#0005# => "0100100000000001",  -- 			LDIH  r0, 0x01   ; r0 := 0x101
      16#0006# => "0101001000000000",  -- 			LD    r2, [r0]   ; 2. Wert in r2
      16#0007# => "0011000000000000",  -- 			XOR   r0, r0, r0
      16#0008# => "0100000000000010",  -- 			LDIL  r0, 0x02
      16#0009# => "0100100000000001",  -- 			LDIH  r0, 0x01   ; r0 := 0x102
      16#000a# => "0011001101101100",  -- 			XOR   r3, r3, r3
      16#000b# => "0011010010010000",  -- 			XOR   r4, r4, r4
      16#000c# => "0100010000000001",  -- 			LDIL  r4, 1
      16#000d# => "0011010110110100",  -- 			XOR   r5, r5, r5
      16#000e# => "0100010100010000",  -- 			LDIL  r5, calc
      16#000f# => "0100110100000000",  -- 			LDIH  r5, calc>>8
      16#0010# => "0000001101100100",  -- calc: 		ADD   r3, r3, r1 ; Addieren, r3 = r3 + r1
      16#0011# => "0000101001010000",  -- 			SUB   r2, r2, r4 ; Subtrahieren, r2 = r2 - r4
      16#0012# => "1001100010101000",  -- 			JNZ   r2, r5
      16#0013# => "0101100000001100",  -- 			ST    [r0], r3   ; Ergebnis speichern
      others => "UUUUUUUUUUUUUUUU"
    );
    
begin
-- Instantiate the Unit Under Test (UUT)
UUT: VISCY_CPU port map (
	clk => clk, reset => reset,
	rd => rd, wr => wr, ready => ready,
	adr => adr, rdata => rdata, wdata => wdata
);
-- Process to simulate the memory behavior...
memory : process
begin
	ready <= '0';
	wait on rd, wr;
		if rd = '1' then
			wait for mem_delay;
			if is_x (adr) then
				rdata <= (others => 'X');
			else
				rdata <= mem_content (to_integer (unsigned (adr)));
			end if;
			ready <= '1';
			wait until rd = '0';
				rdata <= (others => 'X');
			wait for mem_delay;
				ready <= '0';
		elsif wr = '1' then
			wait for mem_delay;
			if not is_x(adr) then
				mem_content (to_integer (unsigned (adr))) <= wdata;
			end if;
			ready <= '1';
			wait until wr = '0';
			wait for mem_delay;
			ready <= '0';
		end if;
end process;

-- Main testbench process...
tb : process
	procedure run_cycle is
	begin
	clk <= '0';
	wait for clk_period / 2;
	clk <= '1';
	wait for clk_period / 2;
	end procedure;
	variable nb_takt: integer :=0;
	begin
	-- SINNVOLLES HAUPTPROGRAMM UEBERLEGEN
		
	reset <= '1';
	run_cycle;
	reset <= '0';
	
	--~ rd <= '1';
	--~ wr <= '0';

	while nb_takt <= 10 loop
		if(rd = '0') then
			nb_takt := nb_takt + 1;
		else
			nb_takt := 0;
		end if;
		run_cycle;
			report "TEST " & integer'image(to_integer(unsigned(adr)));

	end loop;
	wait;
	-- wait forever (stop simulation)
end process;
end;

